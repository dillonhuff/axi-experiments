module top();

   axil_ram #(.DATA_WIDTH(32), .ADDR_WIDTH(5)) ram();
   
endmodule
